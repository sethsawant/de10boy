// converts opcodes into ASCII strings, useful for debugging

module opcode_string (
    input logic [7:0] current_op,
    output reg [24*8-1:0] opcode_str, cb_opcode_str
);
    always@(current_op) begin
        case(current_op)
            8'h00 : opcode_str = "NOP";
            8'h01 : opcode_str = "LD BC d16";
            8'h02 : opcode_str = "LD (BC) A";
            8'h03 : opcode_str = "INC BC";
            8'h04 : opcode_str = "INC B";
            8'h05 : opcode_str = "DEC B";
            8'h06 : opcode_str = "LD B d8";
            8'h07 : opcode_str = "RLCA";
            8'h08 : opcode_str = "LD (a16) SP";
            8'h09 : opcode_str = "ADD HL BC";
            8'h0A : opcode_str = "LD A (BC)";
            8'h0B : opcode_str = "DEC BC";
            8'h0C : opcode_str = "INC C";
            8'h0D : opcode_str = "DEC C";
            8'h0E : opcode_str = "LD C d8";
            8'h0F : opcode_str = "RRCA";
            8'h10 : opcode_str = "STOP";
            8'h11 : opcode_str = "LD DE d16";
            8'h12 : opcode_str = "LD (DE) A";
            8'h13 : opcode_str = "INC DE";
            8'h14 : opcode_str = "INC D";
            8'h15 : opcode_str = "DEC D";
            8'h16 : opcode_str = "LD D d8";
            8'h17 : opcode_str = "RLA";
            8'h18 : opcode_str = "JR r8";
            8'h19 : opcode_str = "ADD HL DE";
            8'h1A : opcode_str = "LD A (DE)";
            8'h1B : opcode_str = "DEC DE";
            8'h1C : opcode_str = "INC E";
            8'h1D : opcode_str = "DEC E";
            8'h1E : opcode_str = "LD E d8";
            8'h1F : opcode_str = "RRA";
            8'h20 : opcode_str = "JR NZ r8";
            8'h21 : opcode_str = "LD HL d16";
            8'h22 : opcode_str = "LD (HL) A";
            8'h23 : opcode_str = "INC HL";
            8'h24 : opcode_str = "INC H";
            8'h25 : opcode_str = "DEC H";
            8'h26 : opcode_str = "LD H d8";
            8'h27 : opcode_str = "DAA";
            8'h28 : opcode_str = "JR Z r8";
            8'h29 : opcode_str = "ADD HL HL";
            8'h2A : opcode_str = "LD A (HL)";
            8'h2B : opcode_str = "DEC HL";
            8'h2C : opcode_str = "INC L";
            8'h2D : opcode_str = "DEC L";
            8'h2E : opcode_str = "LD L d8";
            8'h2F : opcode_str = "CPL";
            8'h30 : opcode_str = "JR NC r8";
            8'h31 : opcode_str = "LD SP d16";
            8'h32 : opcode_str = "LD (HL) A";
            8'h33 : opcode_str = "INC SP";
            8'h34 : opcode_str = "INC (HL)";
            8'h35 : opcode_str = "DEC (HL)";
            8'h36 : opcode_str = "LD (HL) d8";
            8'h37 : opcode_str = "SCF";
            8'h38 : opcode_str = "JR C r8";
            8'h39 : opcode_str = "ADD HL SP";
            8'h3A : opcode_str = "LD A (HL)";
            8'h3B : opcode_str = "DEC SP";
            8'h3C : opcode_str = "INC A";
            8'h3D : opcode_str = "DEC A";
            8'h3E : opcode_str = "LD A d8";
            8'h3F : opcode_str = "CCF";
            8'h40 : opcode_str = "LD B B";
            8'h41 : opcode_str = "LD B C";
            8'h42 : opcode_str = "LD B D";
            8'h43 : opcode_str = "LD B E";
            8'h44 : opcode_str = "LD B H";
            8'h45 : opcode_str = "LD B L";
            8'h46 : opcode_str = "LD B (HL)";
            8'h47 : opcode_str = "LD B A";
            8'h48 : opcode_str = "LD C B";
            8'h49 : opcode_str = "LD C C";
            8'h4A : opcode_str = "LD C D";
            8'h4B : opcode_str = "LD C E";
            8'h4C : opcode_str = "LD C H";
            8'h4D : opcode_str = "LD C L";
            8'h4E : opcode_str = "LD C (HL)";
            8'h4F : opcode_str = "LD C A";
            8'h50 : opcode_str = "LD D B";
            8'h51 : opcode_str = "LD D C";
            8'h52 : opcode_str = "LD D D";
            8'h53 : opcode_str = "LD D E";
            8'h54 : opcode_str = "LD D H";
            8'h55 : opcode_str = "LD D L";
            8'h56 : opcode_str = "LD D (HL)";
            8'h57 : opcode_str = "LD D A";
            8'h58 : opcode_str = "LD E B";
            8'h59 : opcode_str = "LD E C";
            8'h5A : opcode_str = "LD E D";
            8'h5B : opcode_str = "LD E E";
            8'h5C : opcode_str = "LD E H";
            8'h5D : opcode_str = "LD E L";
            8'h5E : opcode_str = "LD E (HL)";
            8'h5F : opcode_str = "LD E A";
            8'h60 : opcode_str = "LD H B";
            8'h61 : opcode_str = "LD H C";
            8'h62 : opcode_str = "LD H D";
            8'h63 : opcode_str = "LD H E";
            8'h64 : opcode_str = "LD H H";
            8'h65 : opcode_str = "LD H L";
            8'h66 : opcode_str = "LD H (HL)";
            8'h67 : opcode_str = "LD H A";
            8'h68 : opcode_str = "LD L B";
            8'h69 : opcode_str = "LD L C";
            8'h6A : opcode_str = "LD L D";
            8'h6B : opcode_str = "LD L E";
            8'h6C : opcode_str = "LD L H";
            8'h6D : opcode_str = "LD L L";
            8'h6E : opcode_str = "LD L (HL)";
            8'h6F : opcode_str = "LD L A";
            8'h70 : opcode_str = "LD (HL) B";
            8'h71 : opcode_str = "LD (HL) C";
            8'h72 : opcode_str = "LD (HL) D";
            8'h73 : opcode_str = "LD (HL) E";
            8'h74 : opcode_str = "LD (HL) H";
            8'h75 : opcode_str = "LD (HL) L";
            8'h76 : opcode_str = "HALT";
            8'h77 : opcode_str = "LD (HL) A";
            8'h78 : opcode_str = "LD A B";
            8'h79 : opcode_str = "LD A C";
            8'h7A : opcode_str = "LD A D";
            8'h7B : opcode_str = "LD A E";
            8'h7C : opcode_str = "LD A H";
            8'h7D : opcode_str = "LD A L";
            8'h7E : opcode_str = "LD A (HL)";
            8'h7F : opcode_str = "LD A A";
            8'h80 : opcode_str = "ADD A B";
            8'h81 : opcode_str = "ADD A C";
            8'h82 : opcode_str = "ADD A D";
            8'h83 : opcode_str = "ADD A E";
            8'h84 : opcode_str = "ADD A H";
            8'h85 : opcode_str = "ADD A L";
            8'h86 : opcode_str = "ADD A (HL)";
            8'h87 : opcode_str = "ADD A A";
            8'h88 : opcode_str = "ADC A B";
            8'h89 : opcode_str = "ADC A C";
            8'h8A : opcode_str = "ADC A D";
            8'h8B : opcode_str = "ADC A E";
            8'h8C : opcode_str = "ADC A H";
            8'h8D : opcode_str = "ADC A L";
            8'h8E : opcode_str = "ADC A (HL)";
            8'h8F : opcode_str = "ADC A A";
            8'h90 : opcode_str = "SUB B";
            8'h91 : opcode_str = "SUB C";
            8'h92 : opcode_str = "SUB D";
            8'h93 : opcode_str = "SUB E";
            8'h94 : opcode_str = "SUB H";
            8'h95 : opcode_str = "SUB L";
            8'h96 : opcode_str = "SUB (HL)";
            8'h97 : opcode_str = "SUB A";
            8'h98 : opcode_str = "SBC A B";
            8'h99 : opcode_str = "SBC A C";
            8'h9A : opcode_str = "SBC A D";
            8'h9B : opcode_str = "SBC A E";
            8'h9C : opcode_str = "SBC A H";
            8'h9D : opcode_str = "SBC A L";
            8'h9E : opcode_str = "SBC A (HL)";
            8'h9F : opcode_str = "SBC A A";
            8'hA0 : opcode_str = "AND B";
            8'hA1 : opcode_str = "AND C";
            8'hA2 : opcode_str = "AND D";
            8'hA3 : opcode_str = "AND E";
            8'hA4 : opcode_str = "AND H";
            8'hA5 : opcode_str = "AND L";
            8'hA6 : opcode_str = "AND (HL)";
            8'hA7 : opcode_str = "AND A";
            8'hA8 : opcode_str = "XOR B";
            8'hA9 : opcode_str = "XOR C";
            8'hAA : opcode_str = "XOR D";
            8'hAB : opcode_str = "XOR E";
            8'hAC : opcode_str = "XOR H";
            8'hAD : opcode_str = "XOR L";
            8'hAE : opcode_str = "XOR (HL)";
            8'hAF : opcode_str = "XOR A";
            8'hB0 : opcode_str = "OR B";
            8'hB1 : opcode_str = "OR C";
            8'hB2 : opcode_str = "OR D";
            8'hB3 : opcode_str = "OR E";
            8'hB4 : opcode_str = "OR H";
            8'hB5 : opcode_str = "OR L";
            8'hB6 : opcode_str = "OR (HL)";
            8'hB7 : opcode_str = "OR A";
            8'hB8 : opcode_str = "CP B";
            8'hB9 : opcode_str = "CP C";
            8'hBA : opcode_str = "CP D";
            8'hBB : opcode_str = "CP E";
            8'hBC : opcode_str = "CP H";
            8'hBD : opcode_str = "CP L";
            8'hBE : opcode_str = "CP (HL)";
            8'hBF : opcode_str = "CP A";
            8'hC0 : opcode_str = "RET NZ";
            8'hC1 : opcode_str = "POP BC";
            8'hC2 : opcode_str = "JP NZ a16";
            8'hC3 : opcode_str = "JP a16";
            8'hC4 : opcode_str = "CALL NZ a16";
            8'hC5 : opcode_str = "PUSH BC";
            8'hC6 : opcode_str = "ADD A d8";
            8'hC7 : opcode_str = "RST 00H";
            8'hC8 : opcode_str = "RET Z";
            8'hC9 : opcode_str = "RET";
            8'hCA : opcode_str = "JP Z a16";
            8'hCB : opcode_str = "PREFIX";
            8'hCC : opcode_str = "CALL Z a16";
            8'hCD : opcode_str = "CALL a16";
            8'hCE : opcode_str = "ADC A d8";
            8'hCF : opcode_str = "RST 08H";
            8'hD0 : opcode_str = "RET NC";
            8'hD1 : opcode_str = "POP DE";
            8'hD2 : opcode_str = "JP NC a16";
            8'hD3 : opcode_str = "ILLEGAL_D3";
            8'hD4 : opcode_str = "CALL NC a16";
            8'hD5 : opcode_str = "PUSH DE";
            8'hD6 : opcode_str = "SUB d8";
            8'hD7 : opcode_str = "RST 10H";
            8'hD8 : opcode_str = "RET C";
            8'hD9 : opcode_str = "RETI";
            8'hDA : opcode_str = "JP C a16";
            8'hDB : opcode_str = "ILLEGAL_DB";
            8'hDC : opcode_str = "CALL C a16";
            8'hDD : opcode_str = "ILLEGAL_DD";
            8'hDE : opcode_str = "SBC A d8";
            8'hDF : opcode_str = "RST 18H";
            8'hE0 : opcode_str = "LDH (a8) A";
            8'hE1 : opcode_str = "POP HL";
            8'hE2 : opcode_str = "LD (C) A";
            8'hE3 : opcode_str = "ILLEGAL_E3";
            8'hE4 : opcode_str = "ILLEGAL_E4";
            8'hE5 : opcode_str = "PUSH HL";
            8'hE6 : opcode_str = "AND d8";
            8'hE7 : opcode_str = "RST 20H";
            8'hE8 : opcode_str = "ADD SP r8";
            8'hE9 : opcode_str = "JP HL";
            8'hEA : opcode_str = "LD (a16) A";
            8'hEB : opcode_str = "ILLEGAL_EB";
            8'hEC : opcode_str = "ILLEGAL_EC";
            8'hED : opcode_str = "ILLEGAL_ED";
            8'hEE : opcode_str = "XOR d8";
            8'hEF : opcode_str = "RST 28H";
            8'hF0 : opcode_str = "LDH A (a8)";
            8'hF1 : opcode_str = "POP AF";
            8'hF2 : opcode_str = "LD A (C)";
            8'hF3 : opcode_str = "DI";
            8'hF4 : opcode_str = "ILLEGAL_F4";
            8'hF5 : opcode_str = "PUSH AF";
            8'hF6 : opcode_str = "OR d8";
            8'hF7 : opcode_str = "RST 30H";
            8'hF8 : opcode_str = "LD HL SP";
            8'hF9 : opcode_str = "LD SP HL";
            8'hFA : opcode_str = "LD A (a16)";
            8'hFB : opcode_str = "EI";
            8'hFC : opcode_str = "ILLEGAL_FC";
            8'hFD : opcode_str = "ILLEGAL_FD";
            8'hFE : opcode_str = "CP d8";
            8'hFF : opcode_str = "RST 38H";
            default : opcode_str = "UKNOWN_OPCODE";
        endcase
    end
    always@(current_op) begin
        case(current_op)
            8'h00 : cb_opcode_str = "RLC B";
            8'h01 : cb_opcode_str = "RLC C";
            8'h02 : cb_opcode_str = "RLC D";
            8'h03 : cb_opcode_str = "RLC E";
            8'h04 : cb_opcode_str = "RLC H";
            8'h05 : cb_opcode_str = "RLC L";
            8'h06 : cb_opcode_str = "RLC (HL)";
            8'h07 : cb_opcode_str = "RLC A";
            8'h08 : cb_opcode_str = "RRC B";
            8'h09 : cb_opcode_str = "RRC C";
            8'h0A : cb_opcode_str = "RRC D";
            8'h0B : cb_opcode_str = "RRC E";
            8'h0C : cb_opcode_str = "RRC H";
            8'h0D : cb_opcode_str = "RRC L";
            8'h0E : cb_opcode_str = "RRC (HL)";
            8'h0F : cb_opcode_str = "RRC A";
            8'h10 : cb_opcode_str = "RL B";
            8'h11 : cb_opcode_str = "RL C";
            8'h12 : cb_opcode_str = "RL D";
            8'h13 : cb_opcode_str = "RL E";
            8'h14 : cb_opcode_str = "RL H";
            8'h15 : cb_opcode_str = "RL L";
            8'h16 : cb_opcode_str = "RL (HL)";
            8'h17 : cb_opcode_str = "RL A";
            8'h18 : cb_opcode_str = "RR B";
            8'h19 : cb_opcode_str = "RR C";
            8'h1A : cb_opcode_str = "RR D";
            8'h1B : cb_opcode_str = "RR E";
            8'h1C : cb_opcode_str = "RR H";
            8'h1D : cb_opcode_str = "RR L";
            8'h1E : cb_opcode_str = "RR (HL)";
            8'h1F : cb_opcode_str = "RR A";
            8'h20 : cb_opcode_str = "SLA B";
            8'h21 : cb_opcode_str = "SLA C";
            8'h22 : cb_opcode_str = "SLA D";
            8'h23 : cb_opcode_str = "SLA E";
            8'h24 : cb_opcode_str = "SLA H";
            8'h25 : cb_opcode_str = "SLA L";
            8'h26 : cb_opcode_str = "SLA (HL)";
            8'h27 : cb_opcode_str = "SLA A";
            8'h28 : cb_opcode_str = "SRA B";
            8'h29 : cb_opcode_str = "SRA C";
            8'h2A : cb_opcode_str = "SRA D";
            8'h2B : cb_opcode_str = "SRA E";
            8'h2C : cb_opcode_str = "SRA H";
            8'h2D : cb_opcode_str = "SRA L";
            8'h2E : cb_opcode_str = "SRA (HL)";
            8'h2F : cb_opcode_str = "SRA A";
            8'h30 : cb_opcode_str = "SWAP B";
            8'h31 : cb_opcode_str = "SWAP C";
            8'h32 : cb_opcode_str = "SWAP D";
            8'h33 : cb_opcode_str = "SWAP E";
            8'h34 : cb_opcode_str = "SWAP H";
            8'h35 : cb_opcode_str = "SWAP L";
            8'h36 : cb_opcode_str = "SWAP (HL)";
            8'h37 : cb_opcode_str = "SWAP A";
            8'h38 : cb_opcode_str = "SRL B";
            8'h39 : cb_opcode_str = "SRL C";
            8'h3A : cb_opcode_str = "SRL D";
            8'h3B : cb_opcode_str = "SRL E";
            8'h3C : cb_opcode_str = "SRL H";
            8'h3D : cb_opcode_str = "SRL L";
            8'h3E : cb_opcode_str = "SRL (HL)";
            8'h3F : cb_opcode_str = "SRL A";
            8'h40 : cb_opcode_str = "BIT 0 B";
            8'h41 : cb_opcode_str = "BIT 0 C";
            8'h42 : cb_opcode_str = "BIT 0 D";
            8'h43 : cb_opcode_str = "BIT 0 E";
            8'h44 : cb_opcode_str = "BIT 0 H";
            8'h45 : cb_opcode_str = "BIT 0 L";
            8'h46 : cb_opcode_str = "BIT 0 (HL)";
            8'h47 : cb_opcode_str = "BIT 0 A";
            8'h48 : cb_opcode_str = "BIT 1 B";
            8'h49 : cb_opcode_str = "BIT 1 C";
            8'h4A : cb_opcode_str = "BIT 1 D";
            8'h4B : cb_opcode_str = "BIT 1 E";
            8'h4C : cb_opcode_str = "BIT 1 H";
            8'h4D : cb_opcode_str = "BIT 1 L";
            8'h4E : cb_opcode_str = "BIT 1 (HL)";
            8'h4F : cb_opcode_str = "BIT 1 A";
            8'h50 : cb_opcode_str = "BIT 2 B";
            8'h51 : cb_opcode_str = "BIT 2 C";
            8'h52 : cb_opcode_str = "BIT 2 D";
            8'h53 : cb_opcode_str = "BIT 2 E";
            8'h54 : cb_opcode_str = "BIT 2 H";
            8'h55 : cb_opcode_str = "BIT 2 L";
            8'h56 : cb_opcode_str = "BIT 2 (HL)";
            8'h57 : cb_opcode_str = "BIT 2 A";
            8'h58 : cb_opcode_str = "BIT 3 B";
            8'h59 : cb_opcode_str = "BIT 3 C";
            8'h5A : cb_opcode_str = "BIT 3 D";
            8'h5B : cb_opcode_str = "BIT 3 E";
            8'h5C : cb_opcode_str = "BIT 3 H";
            8'h5D : cb_opcode_str = "BIT 3 L";
            8'h5E : cb_opcode_str = "BIT 3 (HL)";
            8'h5F : cb_opcode_str = "BIT 3 A";
            8'h60 : cb_opcode_str = "BIT 4 B";
            8'h61 : cb_opcode_str = "BIT 4 C";
            8'h62 : cb_opcode_str = "BIT 4 D";
            8'h63 : cb_opcode_str = "BIT 4 E";
            8'h64 : cb_opcode_str = "BIT 4 H";
            8'h65 : cb_opcode_str = "BIT 4 L";
            8'h66 : cb_opcode_str = "BIT 4 (HL)";
            8'h67 : cb_opcode_str = "BIT 4 A";
            8'h68 : cb_opcode_str = "BIT 5 B";
            8'h69 : cb_opcode_str = "BIT 5 C";
            8'h6A : cb_opcode_str = "BIT 5 D";
            8'h6B : cb_opcode_str = "BIT 5 E";
            8'h6C : cb_opcode_str = "BIT 5 H";
            8'h6D : cb_opcode_str = "BIT 5 L";
            8'h6E : cb_opcode_str = "BIT 5 (HL)";
            8'h6F : cb_opcode_str = "BIT 5 A";
            8'h70 : cb_opcode_str = "BIT 6 B";
            8'h71 : cb_opcode_str = "BIT 6 C";
            8'h72 : cb_opcode_str = "BIT 6 D";
            8'h73 : cb_opcode_str = "BIT 6 E";
            8'h74 : cb_opcode_str = "BIT 6 H";
            8'h75 : cb_opcode_str = "BIT 6 L";
            8'h76 : cb_opcode_str = "BIT 6 (HL)";
            8'h77 : cb_opcode_str = "BIT 6 A";
            8'h78 : cb_opcode_str = "BIT 7 B";
            8'h79 : cb_opcode_str = "BIT 7 C";
            8'h7A : cb_opcode_str = "BIT 7 D";
            8'h7B : cb_opcode_str = "BIT 7 E";
            8'h7C : cb_opcode_str = "BIT 7 H";
            8'h7D : cb_opcode_str = "BIT 7 L";
            8'h7E : cb_opcode_str = "BIT 7 (HL)";
            8'h7F : cb_opcode_str = "BIT 7 A";
            8'h80 : cb_opcode_str = "RES 0 B";
            8'h81 : cb_opcode_str = "RES 0 C";
            8'h82 : cb_opcode_str = "RES 0 D";
            8'h83 : cb_opcode_str = "RES 0 E";
            8'h84 : cb_opcode_str = "RES 0 H";
            8'h85 : cb_opcode_str = "RES 0 L";
            8'h86 : cb_opcode_str = "RES 0 (HL)";
            8'h87 : cb_opcode_str = "RES 0 A";
            8'h88 : cb_opcode_str = "RES 1 B";
            8'h89 : cb_opcode_str = "RES 1 C";
            8'h8A : cb_opcode_str = "RES 1 D";
            8'h8B : cb_opcode_str = "RES 1 E";
            8'h8C : cb_opcode_str = "RES 1 H";
            8'h8D : cb_opcode_str = "RES 1 L";
            8'h8E : cb_opcode_str = "RES 1 (HL)";
            8'h8F : cb_opcode_str = "RES 1 A";
            8'h90 : cb_opcode_str = "RES 2 B";
            8'h91 : cb_opcode_str = "RES 2 C";
            8'h92 : cb_opcode_str = "RES 2 D";
            8'h93 : cb_opcode_str = "RES 2 E";
            8'h94 : cb_opcode_str = "RES 2 H";
            8'h95 : cb_opcode_str = "RES 2 L";
            8'h96 : cb_opcode_str = "RES 2 (HL)";
            8'h97 : cb_opcode_str = "RES 2 A";
            8'h98 : cb_opcode_str = "RES 3 B";
            8'h99 : cb_opcode_str = "RES 3 C";
            8'h9A : cb_opcode_str = "RES 3 D";
            8'h9B : cb_opcode_str = "RES 3 E";
            8'h9C : cb_opcode_str = "RES 3 H";
            8'h9D : cb_opcode_str = "RES 3 L";
            8'h9E : cb_opcode_str = "RES 3 (HL)";
            8'h9F : cb_opcode_str = "RES 3 A";
            8'hA0 : cb_opcode_str = "RES 4 B";
            8'hA1 : cb_opcode_str = "RES 4 C";
            8'hA2 : cb_opcode_str = "RES 4 D";
            8'hA3 : cb_opcode_str = "RES 4 E";
            8'hA4 : cb_opcode_str = "RES 4 H";
            8'hA5 : cb_opcode_str = "RES 4 L";
            8'hA6 : cb_opcode_str = "RES 4 (HL)";
            8'hA7 : cb_opcode_str = "RES 4 A";
            8'hA8 : cb_opcode_str = "RES 5 B";
            8'hA9 : cb_opcode_str = "RES 5 C";
            8'hAA : cb_opcode_str = "RES 5 D";
            8'hAB : cb_opcode_str = "RES 5 E";
            8'hAC : cb_opcode_str = "RES 5 H";
            8'hAD : cb_opcode_str = "RES 5 L";
            8'hAE : cb_opcode_str = "RES 5 (HL)";
            8'hAF : cb_opcode_str = "RES 5 A";
            8'hB0 : cb_opcode_str = "RES 6 B";
            8'hB1 : cb_opcode_str = "RES 6 C";
            8'hB2 : cb_opcode_str = "RES 6 D";
            8'hB3 : cb_opcode_str = "RES 6 E";
            8'hB4 : cb_opcode_str = "RES 6 H";
            8'hB5 : cb_opcode_str = "RES 6 L";
            8'hB6 : cb_opcode_str = "RES 6 (HL)";
            8'hB7 : cb_opcode_str = "RES 6 A";
            8'hB8 : cb_opcode_str = "RES 7 B";
            8'hB9 : cb_opcode_str = "RES 7 C";
            8'hBA : cb_opcode_str = "RES 7 D";
            8'hBB : cb_opcode_str = "RES 7 E";
            8'hBC : cb_opcode_str = "RES 7 H";
            8'hBD : cb_opcode_str = "RES 7 L";
            8'hBE : cb_opcode_str = "RES 7 (HL)";
            8'hBF : cb_opcode_str = "RES 7 A";
            8'hC0 : cb_opcode_str = "SET 0 B";
            8'hC1 : cb_opcode_str = "SET 0 C";
            8'hC2 : cb_opcode_str = "SET 0 D";
            8'hC3 : cb_opcode_str = "SET 0 E";
            8'hC4 : cb_opcode_str = "SET 0 H";
            8'hC5 : cb_opcode_str = "SET 0 L";
            8'hC6 : cb_opcode_str = "SET 0 (HL)";
            8'hC7 : cb_opcode_str = "SET 0 A";
            8'hC8 : cb_opcode_str = "SET 1 B";
            8'hC9 : cb_opcode_str = "SET 1 C";
            8'hCA : cb_opcode_str = "SET 1 D";
            8'hCB : cb_opcode_str = "SET 1 E";
            8'hCC : cb_opcode_str = "SET 1 H";
            8'hCD : cb_opcode_str = "SET 1 L";
            8'hCE : cb_opcode_str = "SET 1 (HL)";
            8'hCF : cb_opcode_str = "SET 1 A";
            8'hD0 : cb_opcode_str = "SET 2 B";
            8'hD1 : cb_opcode_str = "SET 2 C";
            8'hD2 : cb_opcode_str = "SET 2 D";
            8'hD3 : cb_opcode_str = "SET 2 E";
            8'hD4 : cb_opcode_str = "SET 2 H";
            8'hD5 : cb_opcode_str = "SET 2 L";
            8'hD6 : cb_opcode_str = "SET 2 (HL)";
            8'hD7 : cb_opcode_str = "SET 2 A";
            8'hD8 : cb_opcode_str = "SET 3 B";
            8'hD9 : cb_opcode_str = "SET 3 C";
            8'hDA : cb_opcode_str = "SET 3 D";
            8'hDB : cb_opcode_str = "SET 3 E";
            8'hDC : cb_opcode_str = "SET 3 H";
            8'hDD : cb_opcode_str = "SET 3 L";
            8'hDE : cb_opcode_str = "SET 3 (HL)";
            8'hDF : cb_opcode_str = "SET 3 A";
            8'hE0 : cb_opcode_str = "SET 4 B";
            8'hE1 : cb_opcode_str = "SET 4 C";
            8'hE2 : cb_opcode_str = "SET 4 D";
            8'hE3 : cb_opcode_str = "SET 4 E";
            8'hE4 : cb_opcode_str = "SET 4 H";
            8'hE5 : cb_opcode_str = "SET 4 L";
            8'hE6 : cb_opcode_str = "SET 4 (HL)";
            8'hE7 : cb_opcode_str = "SET 4 A";
            8'hE8 : cb_opcode_str = "SET 5 B";
            8'hE9 : cb_opcode_str = "SET 5 C";
            8'hEA : cb_opcode_str = "SET 5 D";
            8'hEB : cb_opcode_str = "SET 5 E";
            8'hEC : cb_opcode_str = "SET 5 H";
            8'hED : cb_opcode_str = "SET 5 L";
            8'hEE : cb_opcode_str = "SET 5 (HL)";
            8'hEF : cb_opcode_str = "SET 5 A";
            8'hF0 : cb_opcode_str = "SET 6 B";
            8'hF1 : cb_opcode_str = "SET 6 C";
            8'hF2 : cb_opcode_str = "SET 6 D";
            8'hF3 : cb_opcode_str = "SET 6 E";
            8'hF4 : cb_opcode_str = "SET 6 H";
            8'hF5 : cb_opcode_str = "SET 6 L";
            8'hF6 : cb_opcode_str = "SET 6 (HL)";
            8'hF7 : cb_opcode_str = "SET 6 A";
            8'hF8 : cb_opcode_str = "SET 7 B";
            8'hF9 : cb_opcode_str = "SET 7 C";
            8'hFA : cb_opcode_str = "SET 7 D";
            8'hFB : cb_opcode_str = "SET 7 E";
            8'hFC : cb_opcode_str = "SET 7 H";
            8'hFD : cb_opcode_str = "SET 7 L";
            8'hFE : cb_opcode_str = "SET 7 (HL)";
            8'hFF : cb_opcode_str = "SET 7 A";
            default : cb_opcode_str = "UKNOWN_OPCODE";
        endcase
    end
endmodule